module snakeoutput(snake);

output [359:0] snake;

assign snake[359:328]=32'd2;
assign snake[295:264]=32'd3;
assign snake[231:200]=32'd1000;

endmodule 